`include "DigitSupply.vh"

module PostLNA
(
  input OuterReceive,
  output InnerReceive,
  input InnerTransmit,
  output OuterTransmit
);


  
endmodule    
