
module GetQDREdge
(
  
