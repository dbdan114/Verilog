`include "DigitSupply.vh"

module OpAmpDO
(
  input V_Plus,
  input input_Plus,
  output output_Plus,
  output output_Minus,
  input input_Minus,
  input V_Minus
);
  tri V_Plus;
  tri input_Plus;
  tri output_Plus;
  tri output_Minus;
  tri input_Minus;
  tri V_Minus;


  
endmodule
