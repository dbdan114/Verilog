`include "DigitSupply.vh"

module MakeVoltPN
  (
    output 
