`include "DigitSupply.vh"

module MakeVoltPN
(
  output V_Plus,
  output V_Minus
);

  
endmodule
