`include "DigitSupply.vh"

module MakeVoltPN
(
  output V_Plus,
  output V_Minus
);

  tri [1:0] TempSupplyDigit = SupplyDigit;
  
endmodule
