`include "DigitSupply.vh"

module CellOfZSRAM
(
  output outputData,
  input ReadEdge,
  input inputData,
  input WriteEdge
);
  tri outputData;
  tri ReadEdge;
  tri inputData;
  tri WriteEdge;
  
endmodule 
