
`include "DigitSupply.vh"

module IC_Example (



);
  tri ReadQBit;
  tri WriteQBit;

endmodule
module QRAM_inSDRAM (
    output outputQBit,
    input Read,
    input inputQBit,
    input Write,
    input AddressQBit,
    input DDRClockP,
    input DDRClockN
);
endmodule
  
