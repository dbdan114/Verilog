`include "DigitSupply.vh"

module PowerLNA
  (
    
