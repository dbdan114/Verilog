`include "DigitSupply.vh"

module CellOfQSRAM
(
  output outputData,
  input ReadEdge,
  input inputData,
  input WriteEdge,
    
  input RefreshEdge
    
);
  tri outputData;
  tri ReadEdge;
  tri inputData;
  tri WriteEdge;
  tri RefreshEdge;

  
  
  _buf MakeInputToSupplyStrength(PreDataToWrite,SupplyDigit,inputData);
endmodule
