module GetQDREdge
(
  output QDREdge,
  input ClockP,
  input ClockN
);
  
endmodule
